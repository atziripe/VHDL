LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RU8 IS
PORT(
		CLK, CLR, CD, CI : IN STD_LOGIC;
		C: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		DATO: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		Q: INOUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE A_RU8 OF RU8 IS
	BEGIN
	
	PROCESS(CLK, CLR)
	BEGIN
		IF(CLR = '0') THEN
			Q <= "000";
		ELSIF(CLK'EVENT AND CLK='1') THEN
			CASE C IS
				WHEN "00" => Q <= DATO;
				WHEN "01" => Q <= Q;
				WHEN "10" =>
							Q <= TO_STDLOGIC(TO_BITVECTOR(Q)) SRL 1)
							Q(7) <= CD;
				WHEN OTHERS =>
							Q <= TO_STDLOGIC(TO_BITVECTOR(Q)) SLL 1)
							Q(7) <= CI;
			END CASE;
		END IF;
	END PROCESS;
END ARCHITECTURE;